module data_memory (
  input  logic        clk,
  input  logic [31:0] address,      // Dirección de memoria
  input  logic [31:0] write_data,   // Datos a escribir
  input  logic        write_enable, // Habilitador de escritura
  input  logic [2:0]  dm_ctrl,      // Control de tamaño y signo
  
  output logic [31:0] read_data,    // Datos leídos
  output logic [31:0] memory_out [0:31] // Salida para debug
);

  // Memoria de datos - 32 palabras (128 bytes)
  logic [31:0] memory [0:31];
  
  // Exponer todas las posiciones para debug
  assign memory_out = memory;

  // Señales intermedias para lectura
  logic [31:0] raw_data;
  logic [7:0]  byte_data;
  logic [15:0] half_data;
  
  // Dirección word-aligned - ASEGURAR QUE ESTÉ EN RANGO
  logic [5:0] word_addr;
  assign word_addr = address[6:2];  // Bits [7:2] para 64 palabras
  // 6:2 → 64 palabras (0-63), 32 palabras en memoria
  // Selección de byte y halfword
  logic [1:0] byte_offset;
  assign byte_offset = address[1:0];
  
  // Lectura de palabra completa - CON PROTECCIÓN DE RANGO
  always_comb begin
    if (word_addr < 64)
      raw_data = memory[word_addr];
    else
      raw_data = 32'hDEADBEEF;  // Valor de debug para direcciones inválidas
  end
  
  // Extracción de byte según offset
  always_comb begin
    case (byte_offset)
      2'b00: byte_data = raw_data[7:0];
      2'b01: byte_data = raw_data[15:8];
      2'b10: byte_data = raw_data[23:16];
      2'b11: byte_data = raw_data[31:24];
      default: byte_data = 8'h00;
    endcase
  end
  
  // Extracción de halfword según offset
  always_comb begin
    case (address[1])
      1'b0: half_data = raw_data[15:0];
      1'b1: half_data = raw_data[31:16];
      default: half_data = 16'h0000;
    endcase
  end
  
  // Control de lectura según dm_ctrl
  always_comb begin
    case (dm_ctrl)
      3'b000: // LB - Load Byte (con signo)
        read_data = {{24{byte_data[7]}}, byte_data};
      
      3'b001: // LH - Load Halfword (con signo)
        read_data = {{16{half_data[15]}}, half_data};
      
      3'b010: // LW - Load Word
        read_data = raw_data;
      
      3'b100: // LBU - Load Byte Unsigned
        read_data = {24'b0, byte_data};
      
      3'b101: // LHU - Load Halfword Unsigned
        read_data = {16'b0, half_data};
      
      default:
        read_data = 32'h00000000;  // Valor por defecto seguro
    endcase
  end
  
  // Escritura síncrona
  always_ff @(posedge clk) begin
    if (write_enable && word_addr < 64) begin
      case (dm_ctrl)
        3'b000: begin // SB - Store Byte
          case (byte_offset)
            2'b00: memory[word_addr][7:0]   <= write_data[7:0];
            2'b01: memory[word_addr][15:8]  <= write_data[7:0];
            2'b10: memory[word_addr][23:16] <= write_data[7:0];
            2'b11: memory[word_addr][31:24] <= write_data[7:0];
          endcase
        end
        
        3'b001: begin // SH - Store Halfword
          case (address[1])
            1'b0: memory[word_addr][15:0]  <= write_data[15:0];
            1'b1: memory[word_addr][31:16] <= write_data[15:0];
          endcase
        end
        
        3'b010: begin // SW - Store Word
          memory[word_addr] <= write_data;
        end
      endcase
    end
  end
  
  // Inicialización con datos de prueba
  initial begin
    // IMPORTANTE: Inicializar TODO el array primero
    for (int i = 0; i < 32; i++) begin
      memory[i] = 32'h00000000;
    end
    
    // Luego establecer valores de prueba
    memory[0]  = 32'h12345678;  // Dirección 0x00
    memory[1]  = 32'hABCDEF00;  // Dirección 0x04
    memory[2]  = 32'h00000064;  // Dirección 0x08 = 100 decimal
    memory[3]  = 32'hFFFFFFFF;  // Dirección 0x0C = -1
    memory[4]  = 32'h000000FF;  // Dirección 0x10 = 255
    memory[5]  = 32'h80000000;  // Dirección 0x14 = número negativo
    
    $display("=== Memoria de datos inicializada ===");
    $display("memory[0] = 0x%h", memory[0]);
    $display("memory[1] = 0x%h", memory[1]);
    $display("memory[2] = 0x%h", memory[2]);
    $display("memory[3] = 0x%h", memory[3]);
  end
  
  // DEBUG: Monitorear lecturas de LW
  always @(posedge clk) begin
    if (!write_enable && dm_ctrl == 3'b010) begin  // LW
      $display("[DEBUG LW] Tiempo=%0t addr=0x%h word_addr=%0d raw_data=0x%h read_data=0x%h", 
               $time, address, word_addr, raw_data, read_data);
    end
  end

endmodule