/*
 * ============================================================
 * Módulo: font_rom
 *
 *   Entrada: addr (11 bits) -> [7 bits ASCII] + [4 bits Fila]
 *   Salida: data (8 bits)   -> Fila de píxeles correspondiente
 * ============================================================
 */

module font_rom (

    input  logic        clk,   
    input  logic [10:0] addr,   // Dirección: Carácter * 16 + Fila
    output logic [7:0]  data    // Datos: 1 = Píxel encendido, 0 = Apagado
	 
);

    logic [7:0] mem [0:2047];
	 
    initial begin
        
        for (int i = 0; i < 2048; i++) begin
            mem[i] = 8'h00;
        end

        // Carácter '&' (ASCII 38)
        mem[38*16 + 3]  = 8'b00110000;
        mem[38*16 + 4]  = 8'b01001000;
        mem[38*16 + 5]  = 8'b01001000;
        mem[38*16 + 6]  = 8'b00110000;
        mem[38*16 + 7]  = 8'b01010100;
        mem[38*16 + 8]  = 8'b01001010;
        mem[38*16 + 9]  = 8'b00110100;

        // Carácter '-' (ASCII 45)
        mem[45*16 + 7]  = 8'b01111100;

        // Carácter ':' (ASCII 58)
        mem[58*16 + 5]  = 8'b00110000;
        mem[58*16 + 9]  = 8'b00110000;

        // Carácter '[' (ASCII 91)
        mem[91*16 + 2]  = 8'b00111100;
        mem[91*16 + 3]  = 8'b00110000;
        mem[91*16 + 4]  = 8'b00110000;
        mem[91*16 + 5]  = 8'b00110000;
        mem[91*16 + 6]  = 8'b00110000;
        mem[91*16 + 7]  = 8'b00110000;
        mem[91*16 + 8]  = 8'b00110000;
        mem[91*16 + 9]  = 8'b00110000;
        mem[91*16 + 10] = 8'b00111100;

        // Carácter ']' (ASCII 93)
        mem[93*16 + 2]  = 8'b00111100;
        mem[93*16 + 3]  = 8'b00001100;
        mem[93*16 + 4]  = 8'b00001100;
        mem[93*16 + 5]  = 8'b00001100;
        mem[93*16 + 6]  = 8'b00001100;
        mem[93*16 + 7]  = 8'b00001100;
        mem[93*16 + 8]  = 8'b00001100;
        mem[93*16 + 9]  = 8'b00001100;
        mem[93*16 + 10] = 8'b00111100;

        // '0' (ASCII 48)
        mem[48*16 + 3]  = 8'b00111100;
        mem[48*16 + 4]  = 8'b01000010;
        mem[48*16 + 5]  = 8'b01000110;
        mem[48*16 + 6]  = 8'b01001010;
        mem[48*16 + 7]  = 8'b01010010;
        mem[48*16 + 8]  = 8'b01100010;
        mem[48*16 + 9]  = 8'b01000010;
        mem[48*16 + 10] = 8'b00111100;

        // '1' (ASCII 49)
        mem[49*16 + 3]  = 8'b00011000;
        mem[49*16 + 4]  = 8'b00111000;
        mem[49*16 + 5]  = 8'b00011000;
        mem[49*16 + 6]  = 8'b00011000;
        mem[49*16 + 7]  = 8'b00011000;
        mem[49*16 + 8]  = 8'b00011000;
        mem[49*16 + 9]  = 8'b00011000;
        mem[49*16 + 10] = 8'b00111100;

        // '2' (ASCII 50)
        mem[50*16 + 3]  = 8'b00111100;
        mem[50*16 + 4]  = 8'b01000010;
        mem[50*16 + 5]  = 8'b00000010;
        mem[50*16 + 6]  = 8'b00000100;
        mem[50*16 + 7]  = 8'b00011000;
        mem[50*16 + 8]  = 8'b00100000;
        mem[50*16 + 9]  = 8'b01000000;
        mem[50*16 + 10] = 8'b01111110;

        // '3' (ASCII 51)
        mem[51*16 + 3]  = 8'b00111100;
        mem[51*16 + 4]  = 8'b01000010;
        mem[51*16 + 5]  = 8'b00000010;
        mem[51*16 + 6]  = 8'b00011100;
        mem[51*16 + 7]  = 8'b00000010;
        mem[51*16 + 8]  = 8'b00000010;
        mem[51*16 + 9]  = 8'b01000010;
        mem[51*16 + 10] = 8'b00111100;

        // '4' (ASCII 52)
        mem[52*16 + 3]  = 8'b00000100;
        mem[52*16 + 4]  = 8'b00001100;
        mem[52*16 + 5]  = 8'b00010100;
        mem[52*16 + 6]  = 8'b00100100;
        mem[52*16 + 7]  = 8'b01000100;
        mem[52*16 + 8]  = 8'b01111110;
        mem[52*16 + 9]  = 8'b00000100;
        mem[52*16 + 10] = 8'b00000100;

        // '5' (ASCII 53)
        mem[53*16 + 3]  = 8'b01111110;
        mem[53*16 + 4]  = 8'b01000000;
        mem[53*16 + 5]  = 8'b01111100;
        mem[53*16 + 6]  = 8'b00000010;
        mem[53*16 + 7]  = 8'b00000010;
        mem[53*16 + 8]  = 8'b00000010;
        mem[53*16 + 9]  = 8'b01000010;
        mem[53*16 + 10] = 8'b00111100;

        // '6' (ASCII 54)
        mem[54*16 + 3]  = 8'b00111100;
        mem[54*16 + 4]  = 8'b01000000;
        mem[54*16 + 5]  = 8'b01000000;
        mem[54*16 + 6]  = 8'b01111100;
        mem[54*16 + 7]  = 8'b01000010;
        mem[54*16 + 8]  = 8'b01000010;
        mem[54*16 + 9]  = 8'b01000010;
        mem[54*16 + 10] = 8'b00111100;

        // '7' (ASCII 55)
        mem[55*16 + 3]  = 8'b01111110;
        mem[55*16 + 4]  = 8'b00000010;
        mem[55*16 + 5]  = 8'b00000100;
        mem[55*16 + 6]  = 8'b00001000;
        mem[55*16 + 7]  = 8'b00010000;
        mem[55*16 + 8]  = 8'b00010000;
        mem[55*16 + 9]  = 8'b00010000;
        mem[55*16 + 10] = 8'b00010000;

        // '8' (ASCII 56)
        mem[56*16 + 3]  = 8'b00111100;
        mem[56*16 + 4]  = 8'b01000010;
        mem[56*16 + 5]  = 8'b01000010;
        mem[56*16 + 6]  = 8'b00111100;
        mem[56*16 + 7]  = 8'b01000010;
        mem[56*16 + 8]  = 8'b01000010;
        mem[56*16 + 9]  = 8'b01000010;
        mem[56*16 + 10] = 8'b00111100;

        // '9' (ASCII 57)
        mem[57*16 + 3]  = 8'b00111100;
        mem[57*16 + 4]  = 8'b01000010;
        mem[57*16 + 5]  = 8'b01000010;
        mem[57*16 + 6]  = 8'b00111110;
        mem[57*16 + 7]  = 8'b00000010;
        mem[57*16 + 8]  = 8'b00000010;
        mem[57*16 + 9]  = 8'b01000010;
        mem[57*16 + 10] = 8'b00111100;

        // 'A' (ASCII 65)
        mem[65*16 + 3]  = 8'b00011000;
        mem[65*16 + 4]  = 8'b00100100;
        mem[65*16 + 5]  = 8'b01000010;
        mem[65*16 + 6]  = 8'b01000010;
        mem[65*16 + 7]  = 8'b01111110;
        mem[65*16 + 8]  = 8'b01000010;
        mem[65*16 + 9]  = 8'b01000010;
        mem[65*16 + 10] = 8'b01000010;

        // 'B' (ASCII 66)
        mem[66*16 + 3]  = 8'b01111100;
        mem[66*16 + 4]  = 8'b01000010;
        mem[66*16 + 5]  = 8'b01000010;
        mem[66*16 + 6]  = 8'b01111100;
        mem[66*16 + 7]  = 8'b01000010;
        mem[66*16 + 8]  = 8'b01000010;
        mem[66*16 + 9]  = 8'b01000010;
        mem[66*16 + 10] = 8'b01111100;

        // 'C' (ASCII 67)
        mem[67*16 + 3]  = 8'b00111100;
        mem[67*16 + 4]  = 8'b01000010;
        mem[67*16 + 5]  = 8'b01000000;
        mem[67*16 + 6]  = 8'b01000000;
        mem[67*16 + 7]  = 8'b01000000;
        mem[67*16 + 8]  = 8'b01000000;
        mem[67*16 + 9]  = 8'b01000010;
        mem[67*16 + 10] = 8'b00111100;

        // 'D' (ASCII 68)
        mem[68*16 + 3]  = 8'b01111000;
        mem[68*16 + 4]  = 8'b01000100;
        mem[68*16 + 5]  = 8'b01000010;
        mem[68*16 + 6]  = 8'b01000010;
        mem[68*16 + 7]  = 8'b01000010;
        mem[68*16 + 8]  = 8'b01000010;
        mem[68*16 + 9]  = 8'b01000100;
        mem[68*16 + 10] = 8'b01111000;

        // 'E' (ASCII 69)
        mem[69*16 + 3]  = 8'b01111110;
        mem[69*16 + 4]  = 8'b01000000;
        mem[69*16 + 5]  = 8'b01000000;
        mem[69*16 + 6]  = 8'b01111100;
        mem[69*16 + 7]  = 8'b01000000;
        mem[69*16 + 8]  = 8'b01000000;
        mem[69*16 + 9]  = 8'b01000000;
        mem[69*16 + 10] = 8'b01111110;

        // 'F' (ASCII 70)
        mem[70*16 + 3]  = 8'b01111110;
        mem[70*16 + 4]  = 8'b01000000;
        mem[70*16 + 5]  = 8'b01000000;
        mem[70*16 + 6]  = 8'b01111100;
        mem[70*16 + 7]  = 8'b01000000;
        mem[70*16 + 8]  = 8'b01000000;
        mem[70*16 + 9]  = 8'b01000000;
        mem[70*16 + 10] = 8'b01000000;

        // 'G' (ASCII 71)
        mem[71*16 + 3]  = 8'b00111100;
        mem[71*16 + 4]  = 8'b01000010;
        mem[71*16 + 5]  = 8'b01000000;
        mem[71*16 + 6]  = 8'b01000000;
        mem[71*16 + 7]  = 8'b01001110;
        mem[71*16 + 8]  = 8'b01000010;
        mem[71*16 + 9]  = 8'b01000010;
        mem[71*16 + 10] = 8'b00111110;

        // 'H' (ASCII 72)
        mem[72*16 + 3]  = 8'b01000010;
        mem[72*16 + 4]  = 8'b01000010;
        mem[72*16 + 5]  = 8'b01000010;
        mem[72*16 + 6]  = 8'b01111110;
        mem[72*16 + 7]  = 8'b01000010;
        mem[72*16 + 8]  = 8'b01000010;
        mem[72*16 + 9]  = 8'b01000010;
        mem[72*16 + 10] = 8'b01000010;

        // 'I' (ASCII 73)
        mem[73*16 + 3]  = 8'b00111000;
        mem[73*16 + 4]  = 8'b00011000;
        mem[73*16 + 5]  = 8'b00011000;
        mem[73*16 + 6]  = 8'b00011000;
        mem[73*16 + 7]  = 8'b00011000;
        mem[73*16 + 8]  = 8'b00011000;
        mem[73*16 + 9]  = 8'b00011000;
        mem[73*16 + 10] = 8'b00111000;

        // 'J' (ASCII 74)
        mem[74*16 + 3]  = 8'b00000110;
        mem[74*16 + 4]  = 8'b00000110;
        mem[74*16 + 5]  = 8'b00000110;
        mem[74*16 + 6]  = 8'b00000110;
        mem[74*16 + 7]  = 8'b00000110;
        mem[74*16 + 8]  = 8'b01000110;
        mem[74*16 + 9]  = 8'b01000110;
        mem[74*16 + 10] = 8'b00111000;

        // 'K' (ASCII 75)
        mem[75*16 + 3]  = 8'b01000010;
        mem[75*16 + 4]  = 8'b01000100;
        mem[75*16 + 5]  = 8'b01001000;
        mem[75*16 + 6]  = 8'b01110000;
        mem[75*16 + 7]  = 8'b01010000;
        mem[75*16 + 8]  = 8'b01001000;
        mem[75*16 + 9]  = 8'b01000100;
        mem[75*16 + 10] = 8'b01000010;

        // 'L' (ASCII 76)
        mem[76*16 + 3]  = 8'b01000000;
        mem[76*16 + 4]  = 8'b01000000;
        mem[76*16 + 5]  = 8'b01000000;
        mem[76*16 + 6]  = 8'b01000000;
        mem[76*16 + 7]  = 8'b01000000;
        mem[76*16 + 8]  = 8'b01000000;
        mem[76*16 + 9]  = 8'b01000000;
        mem[76*16 + 10] = 8'b01111110;

        // 'M' (ASCII 77)
        mem[77*16 + 3]  = 8'b01000010;
        mem[77*16 + 4]  = 8'b01100110;
        mem[77*16 + 5]  = 8'b01011010;
        mem[77*16 + 6]  = 8'b01000010;
        mem[77*16 + 7]  = 8'b01000010;
        mem[77*16 + 8]  = 8'b01000010;
        mem[77*16 + 9]  = 8'b01000010;
        mem[77*16 + 10] = 8'b01000010;

        // 'N' (ASCII 78)
        mem[78*16 + 3]  = 8'b01000010;
        mem[78*16 + 4]  = 8'b01100010;
        mem[78*16 + 5]  = 8'b01010010;
        mem[78*16 + 6]  = 8'b01001010;
        mem[78*16 + 7]  = 8'b01000110;
        mem[78*16 + 8]  = 8'b01000010;
        mem[78*16 + 9]  = 8'b01000010;
        mem[78*16 + 10] = 8'b01000010;

        // 'O' (ASCII 79)
        mem[79*16 + 3]  = 8'b00111100;
        mem[79*16 + 4]  = 8'b01000010;
        mem[79*16 + 5]  = 8'b01000010;
        mem[79*16 + 6]  = 8'b01000010;
        mem[79*16 + 7]  = 8'b01000010;
        mem[79*16 + 8]  = 8'b01000010;
        mem[79*16 + 9]  = 8'b01000010;
        mem[79*16 + 10] = 8'b00111100;

        // 'P' (ASCII 80)
        mem[80*16 + 3]  = 8'b01111100;
        mem[80*16 + 4]  = 8'b01000010;
        mem[80*16 + 5]  = 8'b01000010;
        mem[80*16 + 6]  = 8'b01111100;
        mem[80*16 + 7]  = 8'b01000000;
        mem[80*16 + 8]  = 8'b01000000;
        mem[80*16 + 9]  = 8'b01000000;
        mem[80*16 + 10] = 8'b01000000;

        // 'Q' (ASCII 81)
        mem[81*16 + 3]  = 8'b00111100;
        mem[81*16 + 4]  = 8'b01000010;
        mem[81*16 + 5]  = 8'b01000010;
        mem[81*16 + 6]  = 8'b01000010;
        mem[81*16 + 7]  = 8'b01000010;
        mem[81*16 + 8]  = 8'b01001010;
        mem[81*16 + 9]  = 8'b01000100;
        mem[81*16 + 10] = 8'b00111110;

        // 'R' (ASCII 82)
        mem[82*16 + 3]  = 8'b01111100;
        mem[82*16 + 4]  = 8'b01000010;
        mem[82*16 + 5]  = 8'b01000010;
        mem[82*16 + 6]  = 8'b01111100;
        mem[82*16 + 7]  = 8'b01010000;
        mem[82*16 + 8]  = 8'b01001000;
        mem[82*16 + 9]  = 8'b01000100;
        mem[82*16 + 10] = 8'b01000010;

        // 'S' (ASCII 83)
        mem[83*16 + 3]  = 8'b00111110;
        mem[83*16 + 4]  = 8'b01000000;
        mem[83*16 + 5]  = 8'b01000000;
        mem[83*16 + 6]  = 8'b00111100;
        mem[83*16 + 7]  = 8'b00000010;
        mem[83*16 + 8]  = 8'b00000010;
        mem[83*16 + 9]  = 8'b00000010;
        mem[83*16 + 10] = 8'b01111100;

        // 'T' (ASCII 84)
        mem[84*16 + 3]  = 8'b01111110;
        mem[84*16 + 4]  = 8'b00011000;
        mem[84*16 + 5]  = 8'b00011000;
        mem[84*16 + 6]  = 8'b00011000;
        mem[84*16 + 7]  = 8'b00011000;
        mem[84*16 + 8]  = 8'b00011000;
        mem[84*16 + 9]  = 8'b00011000;
        mem[84*16 + 10] = 8'b00011000;

        // 'U' (ASCII 85)
        mem[85*16 + 3]  = 8'b01000010;
        mem[85*16 + 4]  = 8'b01000010;
        mem[85*16 + 5]  = 8'b01000010;
        mem[85*16 + 6]  = 8'b01000010;
        mem[85*16 + 7]  = 8'b01000010;
        mem[85*16 + 8]  = 8'b01000010;
        mem[85*16 + 9]  = 8'b01000010;
        mem[85*16 + 10] = 8'b00111100;

        // 'V' (ASCII 86)
        mem[86*16 + 3]  = 8'b01000010;
        mem[86*16 + 4]  = 8'b01000010;
        mem[86*16 + 5]  = 8'b01000010;
        mem[86*16 + 6]  = 8'b01000010;
        mem[86*16 + 7]  = 8'b00100100;
        mem[86*16 + 8]  = 8'b00100100;
        mem[86*16 + 9]  = 8'b00011000;
        mem[86*16 + 10] = 8'b00011000;

        // 'W' (ASCII 87)
        mem[87*16 + 3]  = 8'b01000010;
        mem[87*16 + 4]  = 8'b01000010;
        mem[87*16 + 5]  = 8'b01000010;
        mem[87*16 + 6]  = 8'b01000010;
        mem[87*16 + 7]  = 8'b01011010;
        mem[87*16 + 8]  = 8'b01100110;
        mem[87*16 + 9]  = 8'b01000010;

        // 'X' (ASCII 88)
        mem[88*16 + 3]  = 8'b01000010;
        mem[88*16 + 4]  = 8'b00100100;
        mem[88*16 + 5]  = 8'b00100100;
        mem[88*16 + 6]  = 8'b00011000;
        mem[88*16 + 7]  = 8'b00011000;
        mem[88*16 + 8]  = 8'b00100100;
        mem[88*16 + 9]  = 8'b00100100;
        mem[88*16 + 10] = 8'b01000010;

        // 'Y' (ASCII 89)
        mem[89*16 + 3]  = 8'b01000010;
        mem[89*16 + 4]  = 8'b00100100;
        mem[89*16 + 5]  = 8'b00100100;
        mem[89*16 + 6]  = 8'b00011000;
        mem[89*16 + 7]  = 8'b00011000;
        mem[89*16 + 8]  = 8'b00011000;
        mem[89*16 + 9]  = 8'b00011000;
        mem[89*16 + 10] = 8'b00011000;

        // 'Z' (ASCII 90)
        mem[90*16 + 3]  = 8'b01111110;
        mem[90*16 + 4]  = 8'b00000100;
        mem[90*16 + 5]  = 8'b00001000;
        mem[90*16 + 6]  = 8'b00010000;
        mem[90*16 + 7]  = 8'b00100000;
        mem[90*16 + 8]  = 8'b01000000;
        mem[90*16 + 9]  = 8'b01000000;
        mem[90*16 + 10] = 8'b01111110;

        // 'x' (ASCII 120) 
        mem[120*16 + 5]  = 8'b01000010;
        mem[120*16 + 6]  = 8'b00100100;
        mem[120*16 + 7]  = 8'b00011000;
        mem[120*16 + 8]  = 8'b00100100;
        mem[120*16 + 9]  = 8'b01000010;
    end
    
    always_ff @(posedge clk) begin
        data <= mem[addr];
    end

endmodule