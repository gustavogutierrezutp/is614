
module alu (

    input  logic [31:0] A,        // Primer operando
    input  logic [31:0] B,        // Segundo operando
    input  logic [3:0]  ALU_op,   // Selector de operación
    output logic [31:0] ALU_res  // Resultado de la operación     
	 
);

    always_comb begin
	 
        case (ALU_op)
		  
            
            4'b0000: ALU_res = A & B;                          // AND / ANDI
            4'b0001: ALU_res = A | B;                          // OR / ORI
            4'b0011: ALU_res = A ^ B;                          // XOR / XORI

            4'b0010: ALU_res = A + B;                          // ADD / ADDI (Suma)
            4'b0110: ALU_res = A - B;                          // SUB (Resta)

            // Se usan solo los 5 bits menos significativos de B (B[4:0])
            // ya que 2^5 = 32 es el máximo desplazamiento útil.
            4'b0100: ALU_res = A << B[4:0];                    // SLL / SLLI 
            4'b0101: ALU_res = A >> B[4:0];                    // SRL / SRLI 
            4'b0111: ALU_res = $signed(A) >>> B[4:0];          // SRA / SRAI 

            4'b1000: ALU_res = ($signed(A) < $signed(B)) 
                               ? 32'b1 : 32'b0;                // SLT / SLTI (Con signo)
            
            4'b1001: ALU_res = (A < B) ? 32'b1 : 32'b0;        // SLTU / SLTIU (Sin signo)

            // Caso por defecto
            default: ALU_res = 32'b0;
				
        endcase
    end

endmodule