module top_level (
    input  logic [9:0] SW,       // 10 switches de entrada
    input  logic       KEY0,     // botón: 1=unsigned, 0=signed (default)
    output logic [6:0] HEX0,     // nibble bajo
    output logic [6:0] HEX1,     // nibble medio
    output logic [6:0] HEX2,     // nibble medio
    output logic [6:0] HEX3      // nibble alto (incluye signo si aplica)
);

    // ==========================
    // 1) Interpretar el número
    // ==========================
    logic [9:0] unsigned_value;
    logic signed [9:0] signed_value;
    logic signed [10:0] display_value; // un bit más por seguridad

    assign unsigned_value = SW;
    assign signed_value   = SW;

    always_comb begin
        if (KEY0) 
            display_value = unsigned_value; // modo unsigned
        else 
            display_value = signed_value;   // modo signed
    end

    // ==========================
    // 2) Separar en nibbles HEX
    // ==========================
    logic [3:0] nibble0, nibble1, nibble2, nibble3;

    assign nibble0 = display_value[3:0];
    assign nibble1 = display_value[7:4];
    assign nibble2 = {3'b000, display_value[8]};
    assign nibble3 = {3'b000, display_value[9]};

    // ==========================
    // 3) Instanciar decodificadores
    // ==========================
    hex7seg_dec h0 (.bin(nibble0), .seg(HEX0));
    hex7seg_dec h1 (.bin(nibble1), .seg(HEX1));
    hex7seg_dec h2 (.bin(nibble2), .seg(HEX2));
    hex7seg_dec h3 (.bin(nibble3), .seg(HEX3));

endmodule


// ==============================
// Decodificador HEX a 7 segmentos
// ==============================
module hex7seg_dec (
    input  logic [3:0] bin,
    output logic [6:0] seg
);
    always_comb begin
        case (bin)
            4'h0: seg = 7'b1000000; // 0
            4'h1: seg = 7'b1111001; // 1
            4'h2: seg = 7'b0100100; // 2
            4'h3: seg = 7'b0110000; // 3
            4'h4: seg = 7'b0011001; // 4
            4'h5: seg = 7'b0010010; // 5
            4'h6: seg = 7'b0000010; // 6
            4'h7: seg = 7'b1111000; // 7
            4'h8: seg = 7'b0000000; // 8
            4'h9: seg = 7'b0010000; // 9
            4'hA: seg = 7'b0001000; // A
            4'hB: seg = 7'b0000011; // b
            4'hC: seg = 7'b1000110; // C
            4'hD: seg = 7'b0100001; // d
            4'hE: seg = 7'b0000110; // E
            4'hF: seg = 7'b0001110; // F
            default: seg = 7'b1111111; // apagado
        endcase
    end
endmodule
