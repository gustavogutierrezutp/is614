module decoderHEX(

	input [3:0] SW,
	output [6:0] HEX
	
);

assign HEX =  (SW == 4'b0000) ? 7'b1000000 : // 0
              (SW == 4'b0001) ? 7'b1111001 : // 1
              (SW == 4'b0010) ? 7'b0100100 : // 2
              (SW == 4'b0011) ? 7'b0110000 : // 3
              (SW == 4'b0100) ? 7'b0011001 : // 4
              (SW == 4'b0101) ? 7'b0010010 : // 5
              (SW == 4'b0110) ? 7'b0000010 : // 6
              (SW == 4'b0111) ? 7'b1111000 : // 7
              (SW == 4'b1000) ? 7'b0000000 : // 8
              (SW == 4'b1001) ? 7'b0010000 : // 9
              (SW == 4'b1010) ? 7'b0001000 : // A
              (SW == 4'b1011) ? 7'b0000011 : // b
              (SW == 4'b1100) ? 7'b1000110 : // C
              (SW == 4'b1101) ? 7'b0100001 : // d
              (SW == 4'b1110) ? 7'b0000110 : // E
              (SW == 4'b1111) ? 7'b0001110 : // F
                                7'b1111111 ; // Apagado
endmodule