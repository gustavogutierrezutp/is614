module font_rom (
    input  wire        clk,
    input  wire [10:0] addr,
    output reg  [7:0]  data
);

    // ROM embebida - 128 caracteres × 16 filas
    reg [7:0] mem [0:2047];
    
    // Inicialización de la fuente
    initial begin
        integer i;
        
        // Inicializar todo a 0
        for (i = 0; i < 2048; i = i + 1) begin
            mem[i] = 8'h00;
        end
        
        // ========== ESPACIO (32) ==========
        // Ya está en 0
        
        // ========== '&' (38) ==========
        mem[38*16 + 3]  = 8'b00111000;
        mem[38*16 + 4]  = 8'b01101100;
        mem[38*16 + 5]  = 8'b01101100;
        mem[38*16 + 6]  = 8'b00111000;
        mem[38*16 + 7]  = 8'b01110110;
        mem[38*16 + 8]  = 8'b11011100;
        mem[38*16 + 9]  = 8'b11001100;
        mem[38*16 + 10] = 8'b01110110;
        
        // ========== '-' (45) ==========
        mem[45*16 + 7] = 8'b11111110;
        mem[45*16 + 8] = 8'b11111110;
        
        // ========== '0' (48) ==========
        mem[48*16 + 3]  = 8'b00111100;
        mem[48*16 + 4]  = 8'b01100110;
        mem[48*16 + 5]  = 8'b01100110;
        mem[48*16 + 6]  = 8'b01101110;
        mem[48*16 + 7]  = 8'b01110110;
        mem[48*16 + 8]  = 8'b01100110;
        mem[48*16 + 9]  = 8'b01100110;
        mem[48*16 + 10] = 8'b00111100;
        
        // ========== '1' (49) ==========
        mem[49*16 + 3]  = 8'b00011000;
        mem[49*16 + 4]  = 8'b00111000;
        mem[49*16 + 5]  = 8'b00011000;
        mem[49*16 + 6]  = 8'b00011000;
        mem[49*16 + 7]  = 8'b00011000;
        mem[49*16 + 8]  = 8'b00011000;
        mem[49*16 + 9]  = 8'b00011000;
        mem[49*16 + 10] = 8'b01111110;
        
        // ========== '2' (50) ==========
        mem[50*16 + 3]  = 8'b00111100;
        mem[50*16 + 4]  = 8'b01100110;
        mem[50*16 + 5]  = 8'b00000110;
        mem[50*16 + 6]  = 8'b00001100;
        mem[50*16 + 7]  = 8'b00011000;
        mem[50*16 + 8]  = 8'b00110000;
        mem[50*16 + 9]  = 8'b01100000;
        mem[50*16 + 10] = 8'b01111110;
        
        // ========== '3' (51) ==========
        mem[51*16 + 3]  = 8'b00111100;
        mem[51*16 + 4]  = 8'b01100110;
        mem[51*16 + 5]  = 8'b00000110;
        mem[51*16 + 6]  = 8'b00011100;
        mem[51*16 + 7]  = 8'b00000110;
        mem[51*16 + 8]  = 8'b00000110;
        mem[51*16 + 9]  = 8'b01100110;
        mem[51*16 + 10] = 8'b00111100;
        
        // ========== '4' (52) ==========
        mem[52*16 + 3]  = 8'b00001100;
        mem[52*16 + 4]  = 8'b00011100;
        mem[52*16 + 5]  = 8'b00111100;
        mem[52*16 + 6]  = 8'b01101100;
        mem[52*16 + 7]  = 8'b01001100;
        mem[52*16 + 8]  = 8'b01111110;
        mem[52*16 + 9]  = 8'b00001100;
        mem[52*16 + 10] = 8'b00001100;
        
        // ========== '5' (53) ==========
        mem[53*16 + 3]  = 8'b01111110;
        mem[53*16 + 4]  = 8'b01100000;
        mem[53*16 + 5]  = 8'b01111100;
        mem[53*16 + 6]  = 8'b00000110;
        mem[53*16 + 7]  = 8'b00000110;
        mem[53*16 + 8]  = 8'b00000110;
        mem[53*16 + 9]  = 8'b01100110;
        mem[53*16 + 10] = 8'b00111100;
        
        // ========== '6' (54) ==========
        mem[54*16 + 3]  = 8'b00111100;
        mem[54*16 + 4]  = 8'b01100110;
        mem[54*16 + 5]  = 8'b01100000;
        mem[54*16 + 6]  = 8'b01111100;
        mem[54*16 + 7]  = 8'b01100110;
        mem[54*16 + 8]  = 8'b01100110;
        mem[54*16 + 9]  = 8'b01100110;
        mem[54*16 + 10] = 8'b00111100;
        
        // ========== '7' (55) ==========
        mem[55*16 + 3]  = 8'b01111110;
        mem[55*16 + 4]  = 8'b01100110;
        mem[55*16 + 5]  = 8'b00000110;
        mem[55*16 + 6]  = 8'b00001100;
        mem[55*16 + 7]  = 8'b00011000;
        mem[55*16 + 8]  = 8'b00011000;
        mem[55*16 + 9]  = 8'b00011000;
        mem[55*16 + 10] = 8'b00011000;
        
        // ========== '8' (56) ==========
        mem[56*16 + 3]  = 8'b00111100;
        mem[56*16 + 4]  = 8'b01100110;
        mem[56*16 + 5]  = 8'b01100110;
        mem[56*16 + 6]  = 8'b00111100;
        mem[56*16 + 7]  = 8'b01100110;
        mem[56*16 + 8]  = 8'b01100110;
        mem[56*16 + 9]  = 8'b01100110;
        mem[56*16 + 10] = 8'b00111100;
        
        // ========== '9' (57) ==========
        mem[57*16 + 3]  = 8'b00111100;
        mem[57*16 + 4]  = 8'b01100110;
        mem[57*16 + 5]  = 8'b01100110;
        mem[57*16 + 6]  = 8'b01100110;
        mem[57*16 + 7]  = 8'b00111110;
        mem[57*16 + 8]  = 8'b00000110;
        mem[57*16 + 9]  = 8'b01100110;
        mem[57*16 + 10] = 8'b00111100;
        
        // ========== ':' (58) ==========
        mem[58*16 + 5] = 8'b00011000;
        mem[58*16 + 6] = 8'b00011000;
        mem[58*16 + 9] = 8'b00011000;
        mem[58*16 + 10] = 8'b00011000;
        
        // ========== 'A' (65) ==========
        mem[65*16 + 3]  = 8'b00011000;
        mem[65*16 + 4]  = 8'b00111100;
        mem[65*16 + 5]  = 8'b01100110;
        mem[65*16 + 6]  = 8'b01100110;
        mem[65*16 + 7]  = 8'b01111110;
        mem[65*16 + 8]  = 8'b01100110;
        mem[65*16 + 9]  = 8'b01100110;
        mem[65*16 + 10] = 8'b01100110;
        
        // ========== 'B' (66) ==========
        mem[66*16 + 3]  = 8'b01111100;
        mem[66*16 + 4]  = 8'b01100110;
        mem[66*16 + 5]  = 8'b01100110;
        mem[66*16 + 6]  = 8'b01111100;
        mem[66*16 + 7]  = 8'b01100110;
        mem[66*16 + 8]  = 8'b01100110;
        mem[66*16 + 9]  = 8'b01100110;
        mem[66*16 + 10] = 8'b01111100;
        
        // ========== 'C' (67) ==========
        mem[67*16 + 3]  = 8'b00111100;
        mem[67*16 + 4]  = 8'b01100110;
        mem[67*16 + 5]  = 8'b01100000;
        mem[67*16 + 6]  = 8'b01100000;
        mem[67*16 + 7]  = 8'b01100000;
        mem[67*16 + 8]  = 8'b01100000;
        mem[67*16 + 9]  = 8'b01100110;
        mem[67*16 + 10] = 8'b00111100;
        
        // ========== 'D' (68) ==========
        mem[68*16 + 3]  = 8'b01111000;
        mem[68*16 + 4]  = 8'b01101100;
        mem[68*16 + 5]  = 8'b01100110;
        mem[68*16 + 6]  = 8'b01100110;
        mem[68*16 + 7]  = 8'b01100110;
        mem[68*16 + 8]  = 8'b01100110;
        mem[68*16 + 9]  = 8'b01101100;
        mem[68*16 + 10] = 8'b01111000;
        
        // ========== 'E' (69) ==========
        mem[69*16 + 3]  = 8'b01111110;
        mem[69*16 + 4]  = 8'b01100000;
        mem[69*16 + 5]  = 8'b01100000;
        mem[69*16 + 6]  = 8'b01111100;
        mem[69*16 + 7]  = 8'b01100000;
        mem[69*16 + 8]  = 8'b01100000;
        mem[69*16 + 9]  = 8'b01100000;
        mem[69*16 + 10] = 8'b01111110;
        
        // ========== 'F' (70) ==========
        mem[70*16 + 3]  = 8'b01111110;
        mem[70*16 + 4]  = 8'b01100000;
        mem[70*16 + 5]  = 8'b01100000;
        mem[70*16 + 6]  = 8'b01111100;
        mem[70*16 + 7]  = 8'b01100000;
        mem[70*16 + 8]  = 8'b01100000;
        mem[70*16 + 9]  = 8'b01100000;
        mem[70*16 + 10] = 8'b01100000;
        
        // ========== 'G' (71) ==========
        mem[71*16 + 3]  = 8'b00111100;
        mem[71*16 + 4]  = 8'b01100110;
        mem[71*16 + 5]  = 8'b01100000;
        mem[71*16 + 6]  = 8'b01100000;
        mem[71*16 + 7]  = 8'b01101110;
        mem[71*16 + 8]  = 8'b01100110;
        mem[71*16 + 9]  = 8'b01100110;
        mem[71*16 + 10] = 8'b00111100;
        
        // ========== 'H' (72) ==========
        mem[72*16 + 3]  = 8'b01100110;
        mem[72*16 + 4]  = 8'b01100110;
        mem[72*16 + 5]  = 8'b01100110;
        mem[72*16 + 6]  = 8'b01111110;
        mem[72*16 + 7]  = 8'b01100110;
        mem[72*16 + 8]  = 8'b01100110;
        mem[72*16 + 9]  = 8'b01100110;
        mem[72*16 + 10] = 8'b01100110;
        
        // ========== 'I' (73) ==========
        mem[73*16 + 3]  = 8'b00111100;
        mem[73*16 + 4]  = 8'b00011000;
        mem[73*16 + 5]  = 8'b00011000;
        mem[73*16 + 6]  = 8'b00011000;
        mem[73*16 + 7]  = 8'b00011000;
        mem[73*16 + 8]  = 8'b00011000;
        mem[73*16 + 9]  = 8'b00011000;
        mem[73*16 + 10] = 8'b00111100;
        
        // ========== 'J' (74) ==========
        mem[74*16 + 3]  = 8'b00001110;
        mem[74*16 + 4]  = 8'b00000110;
        mem[74*16 + 5]  = 8'b00000110;
        mem[74*16 + 6]  = 8'b00000110;
        mem[74*16 + 7]  = 8'b00000110;
        mem[74*16 + 8]  = 8'b01100110;
        mem[74*16 + 9]  = 8'b01100110;
        mem[74*16 + 10] = 8'b00111100;
        
        // ========== 'K' (75) ==========
        mem[75*16 + 3]  = 8'b01100110;
        mem[75*16 + 4]  = 8'b01101100;
        mem[75*16 + 5]  = 8'b01111000;
        mem[75*16 + 6]  = 8'b01110000;
        mem[75*16 + 7]  = 8'b01111000;
        mem[75*16 + 8]  = 8'b01101100;
        mem[75*16 + 9]  = 8'b01100110;
        mem[75*16 + 10] = 8'b01100110;
        
        // ========== 'L' (76) ==========
        mem[76*16 + 3]  = 8'b01100000;
        mem[76*16 + 4]  = 8'b01100000;
        mem[76*16 + 5]  = 8'b01100000;
        mem[76*16 + 6]  = 8'b01100000;
        mem[76*16 + 7]  = 8'b01100000;
        mem[76*16 + 8]  = 8'b01100000;
        mem[76*16 + 9]  = 8'b01100000;
        mem[76*16 + 10] = 8'b01111110;
        
        // ========== 'M' (77) ==========
        mem[77*16 + 3]  = 8'b01100011;
        mem[77*16 + 4]  = 8'b01110111;
        mem[77*16 + 5]  = 8'b01111111;
        mem[77*16 + 6]  = 8'b01101011;
        mem[77*16 + 7]  = 8'b01100011;
        mem[77*16 + 8]  = 8'b01100011;
        mem[77*16 + 9]  = 8'b01100011;
        mem[77*16 + 10] = 8'b01100011;
        
        // ========== 'N' (78) ==========
        mem[78*16 + 3]  = 8'b01100110;
        mem[78*16 + 4]  = 8'b01110110;
        mem[78*16 + 5]  = 8'b01111110;
        mem[78*16 + 6]  = 8'b01111110;
        mem[78*16 + 7]  = 8'b01101110;
        mem[78*16 + 8]  = 8'b01100110;
        mem[78*16 + 9]  = 8'b01100110;
        mem[78*16 + 10] = 8'b01100110;
        
        // ========== 'O' (79) ==========
        mem[79*16 + 3]  = 8'b00111100;
        mem[79*16 + 4]  = 8'b01100110;
        mem[79*16 + 5]  = 8'b01100110;
        mem[79*16 + 6]  = 8'b01100110;
        mem[79*16 + 7]  = 8'b01100110;
        mem[79*16 + 8]  = 8'b01100110;
        mem[79*16 + 9]  = 8'b01100110;
        mem[79*16 + 10] = 8'b00111100;
        
        // ========== 'P' (80) ==========
        mem[80*16 + 3]  = 8'b01111100;
        mem[80*16 + 4]  = 8'b01100110;
        mem[80*16 + 5]  = 8'b01100110;
        mem[80*16 + 6]  = 8'b01111100;
        mem[80*16 + 7]  = 8'b01100000;
        mem[80*16 + 8]  = 8'b01100000;
        mem[80*16 + 9]  = 8'b01100000;
        mem[80*16 + 10] = 8'b01100000;
        
        // ========== 'Q' (81) ==========
        mem[81*16 + 3]  = 8'b00111100;
        mem[81*16 + 4]  = 8'b01100110;
        mem[81*16 + 5]  = 8'b01100110;
        mem[81*16 + 6]  = 8'b01100110;
        mem[81*16 + 7]  = 8'b01100110;
        mem[81*16 + 8]  = 8'b01101010;
        mem[81*16 + 9]  = 8'b01101100;
        mem[81*16 + 10] = 8'b00110110;
        
        // ========== 'R' (82) ==========
        mem[82*16 + 3]  = 8'b01111100;
        mem[82*16 + 4]  = 8'b01100110;
        mem[82*16 + 5]  = 8'b01100110;
        mem[82*16 + 6]  = 8'b01111100;
        mem[82*16 + 7]  = 8'b01111000;
        mem[82*16 + 8]  = 8'b01101100;
        mem[82*16 + 9]  = 8'b01100110;
        mem[82*16 + 10] = 8'b01100110;
        
        // ========== 'S' (83) ==========
        mem[83*16 + 3]  = 8'b00111100;
        mem[83*16 + 4]  = 8'b01100110;
        mem[83*16 + 5]  = 8'b01100000;
        mem[83*16 + 6]  = 8'b00111100;
        mem[83*16 + 7]  = 8'b00000110;
        mem[83*16 + 8]  = 8'b00000110;
        mem[83*16 + 9]  = 8'b01100110;
        mem[83*16 + 10] = 8'b00111100;
        
        // ========== 'T' (84) ==========
        mem[84*16 + 3]  = 8'b01111110;
        mem[84*16 + 4]  = 8'b00011000;
        mem[84*16 + 5]  = 8'b00011000;
        mem[84*16 + 6]  = 8'b00011000;
        mem[84*16 + 7]  = 8'b00011000;
        mem[84*16 + 8]  = 8'b00011000;
        mem[84*16 + 9]  = 8'b00011000;
        mem[84*16 + 10] = 8'b00011000;
        
        // ========== 'U' (85) ==========
        mem[85*16 + 3]  = 8'b01100110;
        mem[85*16 + 4]  = 8'b01100110;
        mem[85*16 + 5]  = 8'b01100110;
        mem[85*16 + 6]  = 8'b01100110;
        mem[85*16 + 7]  = 8'b01100110;
        mem[85*16 + 8]  = 8'b01100110;
        mem[85*16 + 9]  = 8'b01100110;
        mem[85*16 + 10] = 8'b00111100;
        
        // ========== 'V' (86) ==========
        mem[86*16 + 3]  = 8'b01100110;
        mem[86*16 + 4]  = 8'b01100110;
        mem[86*16 + 5]  = 8'b01100110;
        mem[86*16 + 6]  = 8'b01100110;
        mem[86*16 + 7]  = 8'b01100110;
        mem[86*16 + 8]  = 8'b00111100;
        mem[86*16 + 9]  = 8'b00111100;
        mem[86*16 + 10] = 8'b00011000;
        
        // ========== 'W' (87) ==========
        mem[87*16 + 3]  = 8'b01100011;
        mem[87*16 + 4]  = 8'b01100011;
        mem[87*16 + 5]  = 8'b01100011;
        mem[87*16 + 6]  = 8'b01101011;
        mem[87*16 + 7]  = 8'b01111111;
        mem[87*16 + 8]  = 8'b01110111;
        mem[87*16 + 9]  = 8'b01100011;
        mem[87*16 + 10] = 8'b01100011;
        
        // ========== 'X' (88) ==========
        mem[88*16 + 3]  = 8'b01100110;
        mem[88*16 + 4]  = 8'b01100110;
        mem[88*16 + 5]  = 8'b00111100;
        mem[88*16 + 6]  = 8'b00011000;
        mem[88*16 + 7]  = 8'b00011000;
        mem[88*16 + 8]  = 8'b00111100;
        mem[88*16 + 9]  = 8'b01100110;
        mem[88*16 + 10] = 8'b01100110;
        
        // ========== 'Y' (89) ==========
        mem[89*16 + 3]  = 8'b01100110;
        mem[89*16 + 4]  = 8'b01100110;
        mem[89*16 + 5]  = 8'b01100110;
        mem[89*16 + 6]  = 8'b00111100;
        mem[89*16 + 7]  = 8'b00011000;
        mem[89*16 + 8]  = 8'b00011000;
        mem[89*16 + 9]  = 8'b00011000;
        mem[89*16 + 10] = 8'b00011000;
        
        // ========== 'Z' (90) ==========
        mem[90*16 + 3]  = 8'b01111110;
        mem[90*16 + 4]  = 8'b00000110;
        mem[90*16 + 5]  = 8'b00001100;
        mem[90*16 + 6]  = 8'b00011000;
        mem[90*16 + 7]  = 8'b00110000;
        mem[90*16 + 8]  = 8'b01100000;
        mem[90*16 + 9]  = 8'b01100000;
        mem[90*16 + 10] = 8'b01111110;
        
        // ========== '[' (91) ==========
        mem[91*16 + 2]  = 8'b00111100;
        mem[91*16 + 3]  = 8'b00110000;
        mem[91*16 + 4]  = 8'b00110000;
        mem[91*16 + 5]  = 8'b00110000;
        mem[91*16 + 6]  = 8'b00110000;
        mem[91*16 + 7]  = 8'b00110000;
        mem[91*16 + 8]  = 8'b00110000;
        mem[91*16 + 9]  = 8'b00110000;
        mem[91*16 + 10] = 8'b00111100;
        
        // ========== ']' (93) ==========
        mem[93*16 + 2]  = 8'b00111100;
        mem[93*16 + 3]  = 8'b00001100;
        mem[93*16 + 4]  = 8'b00001100;
        mem[93*16 + 5]  = 8'b00001100;
        mem[93*16 + 6]  = 8'b00001100;
        mem[93*16 + 7]  = 8'b00001100;
        mem[93*16 + 8]  = 8'b00001100;
        mem[93*16 + 9]  = 8'b00001100;
        mem[93*16 + 10] = 8'b00111100;
        
        // ========== 'x' minúscula (120) ==========
        mem[120*16 + 4]  = 8'b01100110;
        mem[120*16 + 5]  = 8'b01100110;
        mem[120*16 + 6]  = 8'b00111100;
        mem[120*16 + 7]  = 8'b00011000;
        mem[120*16 + 8]  = 8'b00111100;
        mem[120*16 + 9]  = 8'b01100110;
        mem[120*16 + 10] = 8'b01100110;
		  
		  // ========== '+' (43) ==========
		  mem[43*16 + 2]  = 8'b00000000;
		  mem[43*16 + 3]  = 8'b00011000;
        mem[43*16 + 4]  = 8'b00011000;
        mem[43*16 + 5]  = 8'b00011000;
        mem[43*16 + 6]  = 8'b01111110;
        mem[43*16 + 7]  = 8'b00011000;
        mem[43*16 + 8]  = 8'b00011000;
        mem[43*16 + 9]  = 8'b00011000;
        mem[43*16 + 10] = 8'b00000000;
    end

    // Lectura síncrona
    always @(posedge clk) begin
        data <= mem[addr];
    end

endmodule