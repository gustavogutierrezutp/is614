module VGA_Display(
	input clock,
	output reg [7:0] vga_red,
	output reg [7:0] vga_green,
	output reg [7:0] vga_blue,
	output vga_hsync,
	output vga_vsync,
	output vga_clock
);

endmodule