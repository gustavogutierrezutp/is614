`timescale 1ns/1ps

module Led1_tb;
    reg [9:0] SW;
    reg       KEY0;
    wire [6:0] HEX0;
    wire [6:0] HEX1;
    wire [6:0] HEX2;
    wire [6:0] HEX3;

    Led1 dut (
        .SW(SW),
        .KEY0(KEY0),   
        .HEX0(HEX0),
        .HEX1(HEX1),
        .HEX2(HEX2),
		  .HEX3(HEX3)
    );

    initial begin
        KEY0 = 1'b1;   // start in UNSIGNED mode
			  SW = 10'b0000000000;			 #10 
			  SW = 10'b0100010001;			 #10 
			  SW = 10'b1000100010;			 #10 
			  SW = 10'b1100110011;			 #10 
			  SW = 10'b1101000100;			 #10 
			  SW = 10'b1101010101;			 #10 
			  SW = 10'b1101100110;			 #10 
			  SW = 10'b1101110111;			 #10 
			  SW = 10'b1110001000;			 #10 
			  SW = 10'b1110011001;			 #10 
			  SW = 10'b1110101010;			 #10 
			  SW = 10'b1110111011;			 #10 
			  SW = 10'b1111001100;			 #10 
			  SW = 10'b1111011101;			 #10 
			  SW = 10'b1111101110;			 #10 
			  SW = 10'b1111111111;			 #10 
			 
        KEY0 = 1'b0;   // start in SIGNED mode
			  SW = 10'b0000000000;			 #10 
			  SW = 10'b0100010001;			 #10 
			  SW = 10'b1000100010;			 #10 
			  SW = 10'b1100110011;			 #10 
			  SW = 10'b1101000100;			 #10 
			  SW = 10'b1101010101;			 #10 
			  SW = 10'b1101100110;			 #10 
			  SW = 10'b1101110111;			 #10 
			  SW = 10'b1110001000;			 #10 
			  SW = 10'b1110011001;			 #10 
			  SW = 10'b1110101010;			 #10 
			  SW = 10'b1110111011;			 #10 
			  SW = 10'b1111001100;			 #10 
			  SW = 10'b1111011101;			 #10 
			  SW = 10'b1111101110;			 #10 
			  SW = 10'b1111111111;			 #10 

        $stop;
    end
endmodule
