module core(
	input wire clk,  //button pulse
	input wire reset,
	output wire [31:0] pc_vga, inst, imm, rs1, rs2, rd, a, b, res, data, out, wrb,
	output [31:0] x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, 
  x29, x30, x31, 
	output [2:0] ctrl, br,
	output [3:0] alu_ctrl
	
);


    // Señales del procesador
    wire [31:0] nextpc, pc, bsum, instruction, mux3a1;
    wire [31:0] rus1, rus2, immext, mux2a1alua, mux2a1alub;
    wire [31:0] alures, datamemory;
    wire [4:0] brop;
    wire [3:0] aluop;
    wire [2:0] immsrc, dmctrl;
    wire [1:0] rudataWrsrc;
    wire aluasrc, alubsrc, ruwr, nextpcsrc, dmwr, clk_vga;

    // Procesador: Componentes internos
    pc program_counter (
        .clk(clk),                   // Reloj
		  .reset(reset),
        .NextPC(nextpc),             // Siguiente PC
        .Pc(pc)                      // PC actual
    );

    sum4 sum (
        .Asum(pc),                   // Valor del PC actual
        .Bsum(bsum)                  // Resultado PC + 4
    );

    instruction_memory instructionmemory (
        .Address(pc),                // Dirección de instrucción
        .Instruction(instruction)    // Instrucción recuperada
    );

    control_unit controlunit (
        .OpCode(instruction[6:0]),
        .Funct3(instruction[14:12]),
        .Funct7(instruction[31:25]),
        .ImmSrc(immsrc),
        .ALUASrc(aluasrc),
        .ALUBSrc(alubsrc),
        .ALUOp(aluop),
        .DMWr(dmwr),
        .DMCtrl(dmctrl),
        .RUDataWrSrc(rudataWrsrc),
        .RUWr(ruwr),
        .BrOp(brop)
    );

    register_unit unidadderegistros (
        .CLK(clk),
		  .reset(reset),
        .rs1(instruction[19:15]),
        .rs2(instruction[24:20]),
        .rd(instruction[11:7]),
        .DataWr(mux3a1),
        .RuWr(ruwr),
        .Rus1(rus1),
        .Rus2(rus2),
		  
		  .x0(x0),
		  .x1(x1),
		  .x2(x2),
		  .x3(x3),
		  .x4(x4),
		  .x5(x5),
		  .x6(x6),
		  .x7(x7),
		  .x8(x8),
		  .x9(x9),
		  .x10(x10),
		  .x11(x11),
		  .x12(x12),
		  .x13(x13),
		  .x14(x14),
		  .x15(x15),
		  .x16(x16),
		  .x17(x17),
		  .x18(x18),
		  .x19(x19),
		  .x20(x20),
		  .x21(x21),
		  .x22(x22),
		  .x23(x23),
		  .x24(x24),
		  .x25(x25),
		  .x26(x26),
		  .x27(x27),
		  .x28(x28),
		  .x29(x29),
		  .x30(x30),
		  .x31(x31)
		  
    );

    imm_generator immgen (
        .Inst(instruction),
        .ImmSrc(immsrc),
        .ImmExt(immext)
    );

    branch_unit branchunit (
        .A(rus1),
        .B(rus2),
        .BrOp(brop),
        .NextPCSrc(nextpcsrc)
    );

    mux_2 mux_2_1_alu_a (
        .A(rus1),
        .B(pc),
        .select(aluasrc),
        .Out(mux2a1alua)
    );

    mux_2 mux_2_1_alu_b (
        .A(rus2),
        .B(immext),
        .select(alubsrc),
        .Out(mux2a1alub)
    );

    alu alu (
        .A(mux2a1alua),
        .B(mux2a1alub),
        .ALUOp(aluop),
        .ALURes(alures)
    );

    mux_2 mux2a1nextpc (
        .A(bsum),
        .B(alures),
        .select(nextpcsrc),
        .Out(nextpc)
    );

    data_memory datamemory_1 (
        .DMWr(dmwr),
        .DMCtrl(dmctrl),
        .Address(alures),
        .DataWr(rus2),
        .DataRd(datamemory)
    );

    mux_3 mux3a1_1 (
        .A(bsum),
        .B(datamemory),
        .C(alures),
        .select(rudataWrsrc),
        .Out(mux3a1)
    );
	 
	 assign inst = instruction;
	 assign pc_vga = pc;	 
	 assign imm = immext;
	 assign rs1 = rus1;
	 assign rs2 = rus2;
	 assign a = mux2a1alua;
	 assign b = mux2a1alub;
	 assign res = alures;
	 assign data = rus2;
	 assign out = datamemory;
	 assign ctrl = dmctrl;
	 assign br = brop;
	 assign wrb = mux3a1;
	 assign alu_ctrl = aluop;

endmodule

